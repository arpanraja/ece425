// ECE 425 MP2: Verilog RTL for Am2901 controller
// Rev 2/17/08

module controller(
	i,					// opcode (add your decoded signals)
	a,b,select_a_hi,select_b_hi,		// decoding of register addresses
	f,c,p,g_lo,p_lo,ovr,z,			// generation of ALU outputs
	y_tri,y_data,oe,			// tristate control of y bus
	ram0,ram3,		// tristate control of RAM shifter
	q0,q3,q0_data,q3_data,			// tristate control of Q shifter
	reg_wr,      //add additiona signals for your design here
	s1L, _s1L, s0L, _s0L, s0ot, _s0ot, inv_s, inv_r, //alu control signals
	s1Q, _s1Q, s0Q, _s0Q,      //Q register input control signals
	s1R, _s1R, s0R, _s0R,
	s1RS, _s1RS, s0RS, _s0RS,
	s1SS, _s1SS, s0SS, _s0SS,
	sY,_sY,
	lo
);

 // define I/O for synthesized control
input [8:0] i;
input [3:0] a, b;
output [15:0] select_a_hi, select_b_hi;
input [3:0] f, c, p;
output g_lo, p_lo, ovr, z;
inout [3:0] y_tri;
input [3:0] y_data;
input oe;
inout ram0, ram3, q0, q3;
input q0_data, q3_data;
output reg_wr;    //define additional I/Os for your design
//alu control signal intialization
output s1L;
output _s1L;
output s0L;
output _s0L;
output s0ot;
output _s0ot;
output inv_s;
output inv_r;
output s1Q, _s1Q, s0Q, _s0Q;
output s1R, _s1R, s0R, _s0R;
output s1RS, _s1RS, s0RS, _s0RS;
output s1SS, _s1SS, s0SS, _s0SS;
output sY,_sY;
output lo;

//alu control signal assignments
assign s1L = ~i[5] & i[4] &i [3];
assign _s1L = ~s1L;
assign s0L = ~i[4];
assign _s0L = ~s0L;
assign s0ot = ~i[5] & (~i[4] | ~i[3]);
assign _s0ot = ~s0ot;
assign inv_r = (i[5] & ~i[4] & ~i[3]) | (~i[5] & i[3]);
assign inv_s = (~i[5] & i[4]) | (i[5] & ~i[4]) | (i[5] & i[3]);
//Q register input control signal assignments
assign s1Q = i[8] & ~i[6];
assign _s1Q = ~s1Q;
assign s0Q = (~i[8] & i[7]) | (i[8] & ~i[7]) | i[6];
assign _s0Q = ~s0Q;
//ram input control signal assignments
assign s1R = ~i[8];
assign _s1R = ~s1R;
assign s0R = ~i[7];
assign _s0R = ~s0R;
//r input control signal assignments
assign s1RS = ~i[2] & ~i[1];
assign _s1RS = ~s1RS;
assign s0RS = (~i[1] & ~i[0]) | ~i[2]; 
assign _s0RS = ~s0RS;

assign s1SS = (~i[2] & ~i[0])|(i[1] & i[0]);
assign _s1SS = ~s1SS;
assign s0SS = (i[1] & ~i[0]) | (~i[2]);
assign _s0SS = ~s0SS;

assign sY = ~i[8] & i[7] & ~i[6];
assign _sY = ~sY;
assign lo = 1'b0;

 // named internal wires carry reusable subexpressions
wire shift_left, shift_right;

 // "assign" statements give us algebraic expressions
assign select_a_hi = 16'h0001 << a;
assign select_b_hi = 16'h0001 << b;
assign shift_left = i[8] & i[7];
assign shift_right = i[8] & ~ i[7];


 // simpler functionality is better implemented directly in logic gates
buf calcg(	g_lo,	~c[3] ); // glitchy with lookahead carry propagation, but shouldn't matter for us :v)
nand calcp(	p_lo,	p[3], p[2], p[1], p[0] );
xor calcovr(	ovr,	c[3], c[2] );
nor calczero(	z,	f[3], f[2], f[1], f[0] );

bufif1 drvy3(	y_tri[3],y_data[3], oe );
bufif1 drvy2(	y_tri[2],y_data[2], oe );
bufif1 drvy1(	y_tri[1],y_data[1], oe );
bufif1 drvy0(	y_tri[0],y_data[0], oe );
bufif1 drvraml( ram3,	f[3], shift_left );
bufif1 drvramr( ram0,	f[0], shift_right );
bufif1 drvqshl( q3,	q3_data, shift_left );
bufif1 drvqshr( q0,	q0_data, shift_right );


 // add your control signals here...
assign reg_wr = i[8] | i[7];
//end

endmodule

